alu
