Arom_inst : Arom PORT MAP (
		address_a	 => address_a_sig,
		address_b	 => address_b_sig,
		clock	 => clock_sig,
		q_a	 => q_a_sig,
		q_b	 => q_b_sig
	);
