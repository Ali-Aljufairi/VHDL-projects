LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

