LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FA IS
	PORT (
		a, b, IN STD_LOGIC;
		c, d : OUT STD_LOGIC);
END ENTITY;

ARCHITECTURE Behavioral OF FA IS
BEGIN

	c <= a XOR b;
	d <= a AND b;

END ARCHITECTURE;