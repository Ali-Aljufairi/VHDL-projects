LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
ENTITY Register_File IS
  PORT (
    Read_Address_1,
    Read_Address_2,
    Write_Address : IN std_logic_vector(2 DOWNTO 0);
    Clk, Rst, WB_enable : IN std_logic;
    write_data : IN std_logic_vector(15 DOWNTO 0);
    Src1_data, Src2_data : OUT std_logic_vector(15 DOWNTO 0)

  );

END ENTITY;

ARCHITECTURE Register_File_Structal OF Register_File IS
  SIGNAL enable : std_logic_vector(7 DOWNTO 0);
  SIGNAL q0, q1, q2, q3, q4, q5, q6, q7 : std_logic_vector(15 DOWNTO 0);

  COMPONENT r_Register IS
    PORT (
      Clk, Rst, enable : IN std_logic;
      d : IN std_logic_vector(15 DOWNTO 0);
      q : OUT std_logic_vector(15 DOWNTO 0)
    );
  END COMPONENT;
BEGIN

  enable <= "00000001" WHEN Write_Address = "000" AND WB_enable = '1' ELSE
    "00000010" WHEN Write_Address = "001" AND WB_enable = '1' ELSE
    "00000100" WHEN Write_Address = "010" AND WB_enable = '1' ELSE
    "00001000" WHEN Write_Address = "011" AND WB_enable = '1' ELSE
    "00010000" WHEN Write_Address = "100" AND WB_enable = '1' ELSE
    "00100000" WHEN Write_Address = "101" AND WB_enable = '1' ELSE
    "01000000" WHEN Write_Address = "110" AND WB_enable = '1' ELSE
    "10000000" WHEN Write_Address = "111" AND WB_enable = '1' ELSE
    "00000000";
  r0 : r_Register PORT MAP(Clk, Rst, enable(0), write_data, q0);
  r1 : r_Register PORT MAP(Clk, Rst, enable(1), write_data, q1);
  r2 : r_Register PORT MAP(Clk, Rst, enable(2), write_data, q2);
  r3 : r_Register PORT MAP(Clk, Rst, enable(3), write_data, q3);
  r4 : r_Register PORT MAP(Clk, Rst, enable(4), write_data, q4);
  r5 : r_Register PORT MAP(Clk, Rst, enable(5), write_data, q5);
  r6 : r_Register PORT MAP(Clk, Rst, enable(6), write_data, q6);
  r7 : r_Register PORT MAP(Clk, Rst, enable(7), write_data, q7);
  Src1_data <= q0 WHEN Read_Address_1 = "000"
    ELSE q1 WHEN Read_Address_1 = "001"
    ELSE q2 WHEN Read_Address_1 = "010"
    ELSE q3 WHEN Read_Address_1 = "011"
    ELSE q4 WHEN Read_Address_1 = "100"
    ELSE q5 WHEN Read_Address_1 = "101"
    ELSE q6 WHEN Read_Address_1 = "110"
    ELSE q7 WHEN Read_Address_1 = "111";
  Src2_data <= q0 WHEN Read_Address_2 = "000"
  
    ELSE q1 WHEN Read_Address_2 = "001"
    ELSE q2 WHEN Read_Address_2 = "010"
    ELSE q3 WHEN Read_Address_2 = "011"
    ELSE q4 WHEN Read_Address_2 = "100"
    ELSE q5 WHEN Read_Address_2 = "101"
    ELSE q6 WHEN Read_Address_2 = "110"
    ELSE q7 WHEN Read_Address_2 = "111";

END ARCHITECTURE;