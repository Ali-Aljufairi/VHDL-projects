LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
ENTITY LOAD_USE_CASE_DETECTOR IS
  PORT (
    EX_MEMR : IN std_logic;
    D_SRC1, D_SRC2, EX_dest : IN std_logic_vector(2 DOWNTO 0);
    LOAD_USE_CASE_OUT : OUT std_logic);
END ENTITY;

ARCHITECTURE LOAD_USE_CASE_DETECTOR_STRUCTURE OF LOAD_USE_CASE_DETECTOR IS
BEGIN

  LOAD_USE_CASE_OUT <= '1' WHEN (EX_MEMR = '1' AND ((EX_dest = D_SRC1) OR (EX_dest = D_SRC2)))
    ELSE
    '0';
END ARCHITECTURE;