library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY COUNTER IS
PORT(
CLK,RST,ENABLE:IN STD_LOGIC;
FINISH_STALLING:OUT STD_LOGIC


);
END ENTITY;

ARCHITECTURE COUNTER_STRUCTRE OF COUNTER IS
SIGNAL COUNT:  integer range 0 to 1;
BEGIN




--PROCESS (CLk) IS
	--BEGIN



	--	IF (rising_edge(CLK) and ENABLE = '1' and RST='0' ) THEN
--COUNT<= COUNT+1;
--if(COUNT=1) then
--Count<='0';
 
--END IF;
--	END PROCESS;

--FINISH_STALLING<='1' when COUNT=1 else
--'0';


END ARCHITECTURE;